/* *****************************************************************************
 * File name: AND8.v
 * Made by: your name here
 * 
 * Description: This file contains the answer to hw3 of class ee271, 2009.
 * ****************************************************************************/


// Put your code here...
module AND8
  (input [7:0] In,
    output Out);


endmodule // AND8

	   
